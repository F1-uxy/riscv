module control_unit (
    input 
);
    
endmodule