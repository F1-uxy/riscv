module programcounter (
    
);
    
endmodule